LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY ALU2 IS
	PORT (A, B :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	      OP :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			neg :OUT STD_LOGIC;
			R1, R2, R3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ALU2;

ARCHITECTURE Behaviour OF ALU2 IS
	SIGNAL result : STD_LOGIC_VECTOR(9 DOWNTO 0);
BEGIN 
	PROCESS(A, B, OP)
	BEGIN
		CASE OP IS
			WHEN "1000000000000000" =>--Increment A by 2
				result <= ("00" & (A + "10"));
				neg <= '0';
			WHEN "0100000000000000" =>--Shift b to the right by 2 units ("concacting 0")
				result<="0000"&B(7)&B(6)&B(5)&B(4)&B(3)&B(2);
				neg <= '0';
			WHEN "0010000000000000" => --Shift A to the right by 4 units ("concacting 1")
				result<="111100"&A(7)&A(6)&A(5)&A(4);
				neg <= '0';
			WHEN "0001000000000000" =>--Find smaller input and output
				IF(A(7 DOWNTO 0)<B(7 DOWNTO 0)) THEN
					result <= "00"&A(7 DOWNTO 0);
				ELSE
					result <= "00"&B(7 DOWNTO 0);
				END IF;
				neg <= '0';
			WHEN "0000100000000000" =>--Rotate A to the right by two bits
				result<="00"&A(1)&A(0)&A(7)&A(6)&A(5)&A(4)&A(3)&A(2);
				neg <= '0';
			WHEN "0000010000000000" =>--Invert bit significance
				result<="00" &B(0)&B(1)&B(2)&B(3)&B(4)&B(5)&B(6)&B(7);
				neg <= '0';
			WHEN "0000001000000000" =>--XOR a and b
				result <= "00" & (A xor B);
				neg <= '0';
			WHEN "0000000100000000" =>--Produce summation of A and B then decrease by 4
				IF (("00" & A) + ("00" & B)<"100")THEN
					result <= not("100"-(("00" & A) + ("00" & B)))+1;
					neg<='1';
				ELSE
					result <= (("00" & A) + ("00" & B)) - "100";
					neg <= '0';
				END IF;
			WHEN "0000000010000000" =>--Output al hig bits
				result <= "1111111111";
				neg <= '0';
			WHEN OTHERS => 
				result <= "1111111111";
		END CASE;
	END PROCESS;
	
	R1 <= "00" & Result(9 DOWNTO 8);
	R2 <= Result(7 DOWNTO 4);
	R3 <= Result(3 DOWNTO 0);
END Behaviour;
	

	
			