library verilog;
use verilog.vl_types.all;
entity Lab6Part2_vlg_vec_tst is
end Lab6Part2_vlg_vec_tst;
